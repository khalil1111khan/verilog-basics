module comparator_2bit(
output G,E,L,
input [1:0]a,b);
assign G = ((a[1]&(~b[1])) | ((~a[1])&a[0]&(~b[1])&(~b[0])) | (a[1]&a[0]&b[1]&(~b[0])));
assign E = (((~a[1])&(~a[0])&(~b[1])&(~b[0])) | ((~a[1])&(a[0])&(~b[1])&(b[0])) | ((a[1])&(~a[0])&(b[1])&(~b[0])) | ((a[1])&(a[0])&(b[1])&(b[0])));
assign L = (((~a[1])&(b[1])) | ((~a[1])&(~a[0])&(~b[1])&(b[0])) | (a[1]&(~a[0])&b[1]&(b[0])));
endmodule
